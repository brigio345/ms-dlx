package specs is
	constant INST_SZ:	integer := 32;
	constant REG_SZ:	integer := 32;
	constant N_REGS:	integer := 32;
end specs;

