package branch_types is
	type branch_t is (
		BRANCH_NO,
		BRANCH_U_R,
		BRANCH_U_A,
		BRANCH_EQ0,
		BRANCH_NE0
	);
end branch_types;

