package source_types is
	type source_t is (
		SOURCE_RF,
		SOURCE_ALU,
		SOURCE_LD
	);
end source_types;

